-------------------------------------------------------------------------------
-- Title       : 
-- Project     : 
-------------------------------------------------------------------------------
-- File        : 
-- Authors     : Joachim Schmidt
-- Company     : Hepia
-- Created     : 
-- Last update : 
-- Platform    : Vivado (synthesis)
-- Standard    : VHDL'08
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2018 Hepia, Geneve
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 01.01.2018   0.0      SCJ 	  Created
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.<PACKAGE_NAME>.all;

